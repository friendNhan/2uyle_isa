module shift_right(// dich trai thanh ghi rs1 di imm bit
  input logic [31:0] rs1,
  input logic [4:0] imm,
  
  output logic [31:0] rd_right
  );
      assign rd_right = 
        (imm==5'b00001)? {1'b0,rs1[31:1]}:
        (imm==5'b00010)? {2'b0,rs1[31:2]}:
        (imm==5'b00011)? {3'b0,rs1[31:3]}:
        (imm==5'b00100)? {4'b0,rs1[31:4]}:
        (imm==5'b00101)? {5'b0,rs1[31:5]}:
        (imm==5'b00110)? {6'b0,rs1[31:6]}:
        (imm==5'b00111)? {7'b0,rs1[31:7]}:
        (imm==5'b01000)? {8'b0,rs1[31:8]}:
        (imm==5'b01001)? {9'b0,rs1[31:9]}:
        (imm==5'b01010)? {10'b0,rs1[31:10]}:
        (imm==5'b01011)? {11'b0,rs1[31:11]}:
        (imm==5'b01100)? {12'b0,rs1[31:12]}:
        (imm==5'b01101)? {13'b0,rs1[31:13]}:
        (imm==5'b01110)? {14'b0,rs1[31:14]}:
        (imm==5'b01111)? {15'b0,rs1[31:15]}:
        (imm==5'b10000)? {16'b0,rs1[31:16]}:
        (imm==5'b10001)? {17'b0,rs1[31:17]}:
        (imm==5'b10010)? {18'b0,rs1[31:18]}:
        (imm==5'b10011)? {19'b0,rs1[31:19]}:
        (imm==5'b10100)? {20'b0,rs1[31:20]}:
        (imm==5'b10101)? {21'b0,rs1[31:21]}:
        (imm==5'b10110)? {22'b0,rs1[31:22]}:
        (imm==5'b10111)? {23'b0,rs1[31:23]}:
        (imm==5'b11000)? {24'b0,rs1[31:24]}:
        (imm==5'b11001)? {25'b0,rs1[31:25]}:
        (imm==5'b11010)? {26'b0,rs1[31:26]}:
        (imm==5'b11011)? {27'b0,rs1[31:27]}:
        (imm==5'b11100)? {28'b0,rs1[31:28]}:           
        (imm==5'b11101)? {29'b0,rs1[31:29]}:
        (imm==5'b11110)? {30'b0,rs1[31:30]}:
        (imm==5'b11111)? {31'b0,rs1[31]}: rs1[31:0];

 endmodule




