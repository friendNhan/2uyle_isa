module shift_left( // dich trai thanh ghi rs1 di imm bit
  input logic [31:0] rs1,
  input logic [4:0] imm,
  
  output logic [31:0] rd_left
  );

    assign rd_left = 
     (imm==5'b00001)? {rs1[30:0],1'b0}:
     (imm==5'b00010)? {rs1[29:0],2'b0}:
     (imm==5'b00011)? {rs1[28:0],3'b0}:
     (imm==5'b00100)? {rs1[27:0],4'b0}:
     (imm==5'b00101)? {rs1[26:0],5'b0}:
     (imm==5'b00110)? {rs1[25:0],6'b0}:
     (imm==5'b00111)? {rs1[24:0],7'b0}:
     (imm==5'b01000)? {rs1[23:0],8'b0}:
     (imm==5'b01001)? {rs1[22:0],9'b0}:
     (imm==5'b01010)? {rs1[21:0],10'b0}:
     (imm==5'b01011)? {rs1[20:0],11'b0}:
     (imm==5'b01100)? {rs1[19:0],12'b0}:
     (imm==5'b01101)? {rs1[18:0],13'b0}:
     (imm==5'b01110)? {rs1[17:0],14'b0}:
     (imm==5'b01111)? {rs1[16:0],15'b0}:
     (imm==5'b10000)? {rs1[15:0],16'b0}:
     (imm==5'b10001)? {rs1[14:0],17'b0}:
     (imm==5'b10010)? {rs1[13:0],18'b0}:
     (imm==5'b10011)? {rs1[12:0],19'b0}:
     (imm==5'b10100)? {rs1[11:0],20'b0}:
     (imm==5'b10101)? {rs1[10:0],21'b0}:
     (imm==5'b10110)? {rs1[9:0],22'b0}:
     (imm==5'b10111)? {rs1[8:0],23'b0}:
     (imm==5'b11000)? {rs1[7:0],24'b0}:
     (imm==5'b11001)? {rs1[6:0],25'b0}:
     (imm==5'b11010)? {rs1[5:0],26'b0}:
     (imm==5'b11011)? {rs1[4:0],27'b0}:
     (imm==5'b11100)? {rs1[3:0],28'b0}:           
     (imm==5'b11101)? {rs1[2:0],29'b0}:
     (imm==5'b11110)? {rs1[1:0],30'b0}:
     (imm==5'b11111)? {rs1[0],31'b0}  : rs1[31:0];	  
 endmodule




