module shift_right_arith(
  input logic [31:0] rs1,
  input logic [4:0] imm,
  
  output logic [31:0] rd_right_arith
  );
      assign rd_right_arith = 
        (imm==5'b00001)? {{rs1[31]},rs1[31:1]}:
        (imm==5'b00010)? {{2{rs1[31]}},rs1[31:2]}:
        (imm==5'b00011)? {{3{rs1[31]}},rs1[31:3]}:
        (imm==5'b00100)? {{4{rs1[31]}},rs1[31:4]}:
        (imm==5'b00101)? {{5{rs1[31]}},rs1[31:5]}:
        (imm==5'b00110)? {{6{rs1[31]}},rs1[31:6]}:
        (imm==5'b00111)? {{7{rs1[31]}},rs1[31:7]}:
        (imm==5'b01000)? {{8{rs1[31]}},rs1[31:8]}:
        (imm==5'b01001)? {{9{rs1[31]}},rs1[31:9]}:
        (imm==5'b01010)? {{10{rs1[31]}},rs1[31:10]}:
        (imm==5'b01011)? {{11{rs1[31]}},rs1[31:11]}:
        (imm==5'b01100)? {{12{rs1[31]}},rs1[31:12]}:
        (imm==5'b01101)? {{13{rs1[31]}},rs1[31:13]}:
        (imm==5'b01110)? {{14{rs1[31]}},rs1[31:14]}:
        (imm==5'b01111)? {{15{rs1[31]}},rs1[31:15]}:
        (imm==5'b10000)? {{16{rs1[31]}},rs1[31:16]}:
        (imm==5'b10001)? {{17{rs1[31]}},rs1[31:17]}:
        (imm==5'b10010)? {{18{rs1[31]}},rs1[31:18]}:
        (imm==5'b10011)? {{19{rs1[31]}},rs1[31:19]}:
        (imm==5'b10100)? {{20{rs1[31]}},rs1[31:20]}:
        (imm==5'b10101)? {{21{rs1[31]}},rs1[31:21]}:
        (imm==5'b10110)? {{22{rs1[31]}},rs1[31:22]}:
        (imm==5'b10111)? {{23{rs1[31]}},rs1[31:23]}:
        (imm==5'b11000)? {{24{rs1[31]}},rs1[31:24]}:
        (imm==5'b11001)? {{25{rs1[31]}},rs1[31:25]}:
        (imm==5'b11010)? {{26{rs1[31]}},rs1[31:26]}:
        (imm==5'b11011)? {{27{rs1[31]}},rs1[31:27]}:
        (imm==5'b11100)? {{28{rs1[31]}},rs1[31:28]}:           
        (imm==5'b11101)? {{29{rs1[31]}},rs1[31:29]}:
        (imm==5'b11110)? {{30{rs1[31]}},rs1[31:30]}:
        (imm==5'b11111)? {32{rs1[31]}}					: rs1[31:0];

 endmodule




